//---------------------------------------------------------------------
// Jason Wilden 2025
//---------------------------------------------------------------------
`default_nettype none

module midi_parser (                              // MIDI parser
  
);



endmodule