//---------------------------------------------------------------------
// Jason Wilden 2025
//---------------------------------------------------------------------
`default_nettype none

module midi_parser (                              // MIDI parser
  input var logic i_clk,
  input var logic i_reset_n
);



endmodule